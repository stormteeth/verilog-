module shift_reg(reg_out,reg_in,clock)
output[3:0]reg_out;
intput[3:0]reg_in;
input clock;
endmodule